module clk_metadata_adapter_v1_0_0 
( 
	input clk_in,
	output clk_out
);

    assign clk_out=clk_in;

endmodule


